module Cars_Movement(
);
endmodule